`include "CONSTANTS.v"
module ROM_Lookup(input [4:0] index ,
    input [1:0] mode, //LINEAR = 00 , CIRCULAR = 10, HYPERBOLIC = 11
    output [31:0] module_output);

  
    wire [31:0] atan_table [0:31];
    wire [31:0] atanh_table [0:31];
    wire [31:0] lin_table [0:31];

//00010000000000000000000000000000 45 deg
//00110000000000000000000000000000 135 deg
//01010000000000000000000000000000 225 deg
//01110000000000000000000000000000 315 deg

    assign atan_table[0] 	= 32'b00010000000000000000000000000000;
    assign atan_table[1] 	= 32'b00001001011100100000001010001111;
    assign atan_table[2] 	= 32'b00000100111111011001110000101110;
    assign atan_table[3] 	= 32'b00000010100010001000100011101010;
    assign atan_table[4] 	= 32'b00000001010001011000011010100010;
    assign atan_table[5] 	= 32'b00000000101000101110101111110001;
    assign atan_table[6] 	= 32'b00000000010100010111101100001111;
    assign atan_table[7] 	= 32'b00000000001010001011111000101011;
    assign atan_table[8] 	= 32'b00000000000101000101111100101010;
    assign atan_table[9] 	= 32'b00000000000010100010111110010111;
    assign atan_table[10] 	= 32'b00000000000001010001011111001100;
    assign atan_table[11] 	= 32'b00000000000000101000101111100110;
    assign atan_table[12] 	= 32'b00000000000000010100010111110011;
    assign atan_table[13] 	= 32'b00000000000000001010001011111010;
    assign atan_table[14] 	= 32'b00000000000000000101000101111101;
    assign atan_table[15] 	= 32'b00000000000000000010100010111110;
    assign atan_table[16] 	= 32'b00000000000000000001010001011111;
    assign atan_table[17] 	= 32'b00000000000000000000101000110000;
    assign atan_table[18] 	= 32'b00000000000000000000010100011000;
    assign atan_table[19] 	= 32'b00000000000000000000001010001100;
    assign atan_table[20] 	= 32'b00000000000000000000000101000110;
    assign atan_table[21] 	= 32'b00000000000000000000000010100011;
    assign atan_table[22] 	= 32'b00000000000000000000000001010001;
    assign atan_table[23] 	= 32'b00000000000000000000000000101001;
    assign atan_table[24] 	= 32'b00000000000000000000000000010100;
    assign atan_table[25] 	= 32'b00000000000000000000000000001010;
    assign atan_table[26] 	= 32'b00000000000000000000000000000101;
    assign atan_table[27] 	= 32'b00000000000000000000000000000011;
    assign atan_table[28] 	= 32'b00000000000000000000000000000001;
    assign atan_table[29] 	= 32'b00000000000000000000000000000001;
    assign atan_table[30] 	= 32'b00000000000000000000000000000000;
    assign atan_table[31] 	= 32'b00000000000000000000000000000000;

    assign atanh_table[0] 	= 32'b01000110010011111010100111101011; //dont now what is this exactly
    assign atanh_table[1] 	= 32'b01000110010011111010100111101011;
    assign atanh_table[2] 	= 32'b00100000101100010101110111110101;
    assign atanh_table[3] 	= 32'b00010000000101011000100100011101;
    assign atanh_table[4] 	= 32'b00001000000000101010110001000101;
    assign atanh_table[5] 	= 32'b00000100000000000101010101100010;
    assign atanh_table[6] 	= 32'b00000010000000000000101010101011;
    assign atanh_table[7] 	= 32'b00000001000000000000000101010101;
    assign atanh_table[8] 	= 32'b00000000100000000000000000101011;
    assign atanh_table[9] 	= 32'b00000000010000000000000000000101;
    assign atanh_table[10] 	= 32'b00000000001000000000000000000001;
    assign atanh_table[11] 	= 32'b00000000000100000000000000000000;
    assign atanh_table[12] 	= 32'b00000000000010000000000000000000;
    assign atanh_table[13] 	= 32'b00000000000001000000000000000000;
    assign atanh_table[14] 	= 32'b00000000000000100000000000000000;
    assign atanh_table[15] 	= 32'b00000000000000010000000000000000;
    assign atanh_table[16] 	= 32'b00000000000000001000000000000000;
    assign atanh_table[17] 	= 32'b00000000000000000100000000000000;
    assign atanh_table[18] 	= 32'b00000000000000000010000000000000;
    assign atanh_table[19] 	= 32'b00000000000000000001000000000000;
    assign atanh_table[20] 	= 32'b00000000000000000000100000000000;
    assign atanh_table[21] 	= 32'b00000000000000000000010000000000;
    assign atanh_table[22] 	= 32'b00000000000000000000001000000000;
    assign atanh_table[23] 	= 32'b00000000000000000000000100000000;
    assign atanh_table[24] 	= 32'b00000000000000000000000010000000;
    assign atanh_table[25] 	= 32'b00000000000000000000000001000000;
    assign atanh_table[26] 	= 32'b00000000000000000000000000100000;
    assign atanh_table[27] 	= 32'b00000000000000000000000000010000;
    assign atanh_table[28] 	= 32'b00000000000000000000000000001000;
    assign atanh_table[29] 	= 32'b00000000000000000000000000000100;
    assign atanh_table[30] 	= 32'b00000000000000000000000000000010;
    assign atanh_table[31] 	= 32'b00000000000000000000000000000001;


    assign lin_table[0] 	= 32'b10000000000000000000000000000000;
    assign lin_table[1] 	= 32'b01000000000000000000000000000000;
    assign lin_table[2] 	= 32'b00100000000000000000000000000000;
    assign lin_table[3] 	= 32'b00010000000000000000000000000000;
    assign lin_table[4] 	= 32'b00001000000000000000000000000000;
    assign lin_table[5] 	= 32'b00000100000000000000000000000000;
    assign lin_table[6] 	= 32'b00000010000000000000000000000000;
    assign lin_table[7] 	= 32'b00000001000000000000000000000000;
    assign lin_table[8] 	= 32'b00000000100000000000000000000000;
    assign lin_table[9] 	= 32'b00000000010000000000000000000000;
    assign lin_table[10] 	= 32'b00000000001000000000000000000000;
    assign lin_table[11] 	= 32'b00000000000100000000000000000000;
    assign lin_table[12] 	= 32'b00000000000010000000000000000000;
    assign lin_table[13] 	= 32'b00000000000001000000000000000000;
    assign lin_table[14] 	= 32'b00000000000000100000000000000000;
    assign lin_table[15] 	= 32'b00000000000000010000000000000000;
    assign lin_table[16] 	= 32'b00000000000000001000000000000000;
    assign lin_table[17] 	= 32'b00000000000000000100000000000000;
    assign lin_table[18] 	= 32'b00000000000000000010000000000000;
    assign lin_table[19] 	= 32'b00000000000000000001000000000000;
    assign lin_table[20] 	= 32'b00000000000000000000100000000000;
    assign lin_table[21] 	= 32'b00000000000000000000010000000000;
    assign lin_table[22] 	= 32'b00000000000000000000001000000000;
    assign lin_table[23] 	= 32'b00000000000000000000000100000000;
    assign lin_table[24] 	= 32'b00000000000000000000000010000000;
    assign lin_table[25] 	= 32'b00000000000000000000000001000000;
    assign lin_table[26] 	= 32'b00000000000000000000000000100000;
    assign lin_table[27] 	= 32'b00000000000000000000000000010000;
    assign lin_table[28] 	= 32'b00000000000000000000000000001000;
    assign lin_table[29] 	= 32'b00000000000000000000000000000100;
    assign lin_table[30] 	= 32'b00000000000000000000000000000010;
    assign lin_table[31] 	= 32'b00000000000000000000000000000001;






    assign module_output = (mode == `CIRCULAR)? atan_table[index] : ((mode == `HYPERBOLIC)? atanh_table[index] : lin_table[index]);

endmodule

